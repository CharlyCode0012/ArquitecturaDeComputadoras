//Lozano Carlos Daniel 224003566
//1.- definir modulo y uss i/O
module _and (input A, input B, output C);
//2.- declarar señales/elementos internos

/*3.-comportamiento/implementacion del modulo 
(asiganciones, instancias, conexiones)
*/
assign C = A & B;
//4.- Compilar y si ya esta la palomita verde vamos a library
//5.- 

endmodule
