module CicloFetch();

endmodule