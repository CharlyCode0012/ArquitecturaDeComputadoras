module PC();
endmodule