module();
	
endmodule;