//Lozano Carlos Daniel 224003566
//https://github.com/CharlyCode0012/ArquitecturaDeComputadoras.git

module _nand (input A, input B, output C);

assign C = ~(A & B);


endmodule
