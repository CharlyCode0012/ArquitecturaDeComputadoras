module Sum(op1, op2, result);
input op1, op2;
output result;

assign result = op1 + op2;
endmodule