module MemInstrucciones(input [31:0] DirIn, output[31:0]Instr);
    reg [31:0] Mem [0:255];

    
endmodule