//Lozano Carlos Daniel 224003566
//https://github.com/CharlyCode0012/ArquitecturaDeComputadoras.git

module _or (input A, input B, output C);

assign C = A | B;


endmodule
