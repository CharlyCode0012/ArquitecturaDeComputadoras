module fullSum(input [3:0]A, [3:0]B, [3:0]C, output [3:0]C);


endmodule