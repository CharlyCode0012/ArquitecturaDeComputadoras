//Lozano Carlos Daniel 224003566
//https://github.com/CharlyCode0012/ArquitecturaDeComputadoras.git

module _not (input A, output B);

assign B = ~A;


endmodule
