//Lozano Carlos Daniel 224003566
//https://github.com/CharlyCode0012/ArquitecturaDeComputadoras.git

module _yes (input A, output B);

assign B = A;


endmodule
